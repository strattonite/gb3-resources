

`include "../include/rv32i-defines.v"
`include "../include/sail-core-defines.v"



/*
 *	Description:
 *
 *		This module implements the ALU for the RV32I.
 */



/*
 *	Not all instructions are fed to the ALU. As a result, the ALUctl
 *	field is only unique across the instructions that are actually
 *	fed to the ALU.
 */
module alu(ALUctl, A, B, ALUOut, Branch_Enable, alu_enable);
	input [6:0]		ALUctl;
	input [31:0]		A;
	input [31:0]		B;
	input 			alu_enable;
	output reg [31:0]	ALUOut;
	output reg		Branch_Enable;

	wire [31:0] sum;
	wire [31:0] sub;

    dsp_add add_inst(
        .a_in(A),
        .b_in(B),
        .sum(sum),
    );

    dsp_sub sub_inst(
        .a_in(A),
        .b_in(B),
        .sub(sub),
    );

	/*
	 *	This uses Yosys's support for nonzero initial values:
	 *
	 *		https://github.com/YosysHQ/yosys/commit/0793f1b196df536975a044a4ce53025c81d00c7f
	 *
	 *	Rather than using this simulation construct (`initial`),
	 *	the design should instead use a reset signal going to
	 *	modules in the design.
	 */
	initial begin
		ALUOut = 32'b0;
		Branch_Enable = 1'b0;
	end

	always @(ALUctl, A, B) begin
		if(alu_enable) begin
			case (ALUctl[3:0])
				/*
				*	AND (the fields also match ANDI and LUI)
				*/
				`kSAIL_MICROARCHITECTURE_ALUCTL_3to0_AND:	ALUOut = A & B;

				/*
				*	OR (the fields also match ORI)
				*/
				`kSAIL_MICROARCHITECTURE_ALUCTL_3to0_OR:	ALUOut = A | B;

				/*
				*	ADD (the fields also match AUIPC, all loads, all stores, and ADDI)
				*/
				`kSAIL_MICROARCHITECTURE_ALUCTL_3to0_ADD:	ALUOut = sum;

				/*
				*	SUBTRACT (the fields also matches all branches)
				*/
				`kSAIL_MICROARCHITECTURE_ALUCTL_3to0_SUB:	ALUOut = sub;

				/*
				*	SLT (the fields also matches all the other SLT variants)
				*/
				`kSAIL_MICROARCHITECTURE_ALUCTL_3to0_SLT:	ALUOut = $signed(A) < $signed(B) ? 32'b1 : 32'b0;

				/*
				*	SRL (the fields also matches the other SRL variants)
				*/
				`kSAIL_MICROARCHITECTURE_ALUCTL_3to0_SRL:	ALUOut = A >> B[4:0];

				/*
				*	SRA (the fields also matches the other SRA variants)
				*/
				`kSAIL_MICROARCHITECTURE_ALUCTL_3to0_SRA:	ALUOut = $signed(A) >>> B[4:0];

				/*
				*	SLL (the fields also match the other SLL variants)
				*/
				`kSAIL_MICROARCHITECTURE_ALUCTL_3to0_SLL:	ALUOut = A << B[4:0];

				/*
				*	XOR (the fields also match other XOR variants)
				*/
				`kSAIL_MICROARCHITECTURE_ALUCTL_3to0_XOR:	ALUOut = A ^ B;

				/*
				*	CSRRW  only
				*/
				`kSAIL_MICROARCHITECTURE_ALUCTL_3to0_CSRRW:	ALUOut = A;

				/*
				*	CSRRS only
				*/
				`kSAIL_MICROARCHITECTURE_ALUCTL_3to0_CSRRS:	ALUOut = A | B;

				/*
				*	CSRRC only
				*/
				`kSAIL_MICROARCHITECTURE_ALUCTL_3to0_CSRRC:	ALUOut = (~A) & B;

				/*
				*	Should never happen.
				*/
				default:					ALUOut = 0;
			endcase
		end
		else begin
			ALUOut = 32'b0; // Set to a constant value when alu_enable = 0
		end

	always @(ALUctl, ALUOut, A, B) begin
		case (ALUctl[6:4])
			`kSAIL_MICROARCHITECTURE_ALUCTL_6to4_BEQ:	Branch_Enable = (ALUOut == 0);
			`kSAIL_MICROARCHITECTURE_ALUCTL_6to4_BNE:	Branch_Enable = !(ALUOut == 0);
			`kSAIL_MICROARCHITECTURE_ALUCTL_6to4_BLT:	Branch_Enable = ($signed(A) < $signed(B));
			`kSAIL_MICROARCHITECTURE_ALUCTL_6to4_BGE:	Branch_Enable = ($signed(A) >= $signed(B));
			`kSAIL_MICROARCHITECTURE_ALUCTL_6to4_BLTU:	Branch_Enable = ($unsigned(A) < $unsigned(B));
			`kSAIL_MICROARCHITECTURE_ALUCTL_6to4_BGEU:	Branch_Enable = ($unsigned(A) >= $unsigned(B));

			default:					Branch_Enable = 1'b0;
		endcase
	end
endmodule
